module pl_ddr_top
(

);
endmodule